
library ieee;
use ieee.std_logic_1164.all;

library work;
use work.bus_pkg.all;

package imotor_module_pkg is

   type parity_type is (None, Even, Odd);
   
   -- components here!

end imotor_module_pkg;
