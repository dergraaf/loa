../../../../roboter/2012_captain/software/projects/beacon_system/beacon/fpga_memory_map.vhd