../../../../roboter/2012_captain/software/projects/beacon_system/beacon_test/fpga_memory_map.vhd