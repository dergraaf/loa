../../../../beacon/big/generated/fpga_memory_map.vhd